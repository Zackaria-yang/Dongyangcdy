//****************************************Copyright (c)***********************************//
//ԭ�Ӹ����߽�ѧƽ̨��www.yuanzige.com
//����֧�֣�www.openedv.com
//�Ա����̣�http://openedv.taobao.com
//��ע΢�Ź���ƽ̨΢�źţ�"����ԭ��"����ѻ�ȡZYNQ & FPGA & STM32 & LINUX���ϡ�
//��Ȩ���У�����ؾ���
//Copyright(C) ����ԭ�� 2018-2028
//All rights reserved
//----------------------------------------------------------------------------------------
// File name:           scale_top
// Last modified Date:  2020/09/04 9:19:08
// Last Version:        V1.0
// Descriptions:        ͼ�����Ŷ����װģ��	
//                      
//----------------------------------------------------------------------------------------
// Created by:          ����ԭ��
// Created date:        2020/09/04 9:19:08
// Version:             V1.0
// Descriptions:        The original version
//
//----------------------------------------------------------------------------------------
//****************************************************************************************//

module vip_scale(
	input 			pixel_clk,     //ԭʼ����ʱ��
	input 			sram_clk,      //���ź�����ʱ��
	input           sys_rst_n,     //��λ�ź�	
	input 			hs,            //���ź�
	input 			vs,            //���ź�
	input 			de,            //����ʹ���ź� 
	input	[11:0]  s_width,       //����ǰ���
	input	[11:0]  s_height,      //����ǰ�߶�
	input	[11:0]  t_width,       //���ź���
	input	[11:0]  t_height,	   //���ź�߶� 
	input   [15:0]  h_scale_k,     //����������
	input   [15:0]  v_scale_k,	   //����������	
	input	[15:0]	pixel_data,    //����ǰ����
	output	[15:0]  sram_data_out, //���ź�����
	output  		data_valid     //���ź�������Ч�ź�
    );

//wire define    
wire [15:0] sram_data_out;  //���ź��RGB����
wire [7:0]  data_out_r;     //���ź�ĺ�ɫ����
wire [7:0]  data_out_g;     //���ź����ɫ����
wire [7:0]  data_out_b;     //���ź����ɫ����
wire        data_valid;     //���ź�������Ч�ź�

//*****************************************************
//**                    main code
//*****************************************************

//�����ź������ƴ��16bit�������    
assign  sram_data_out = data_valid ? {data_out_r[7:3],data_out_g[7:2],data_out_b[7:3]} : 16'b0; 
assign  fifo_rden = ~fifo_empty_r && ~fifo_empty_g && ~fifo_empty_b;    

//��ɫ��������ģ��    
 vin_scale_down u_vin_scale_down_r(
	.pixel_clk          (pixel_clk),
	.sram_clk           (sram_clk),
	.sys_rst_n          (sys_rst_n),
	.hs                 (hs),
	.vs                 (vs),
	.de                 (de),
    .s_width            (s_width),
    .s_height           (s_height),
    .t_width            (t_width),
    .t_height           (t_height),
	.h_scale_k          (h_scale_k),
	.v_scale_k          (v_scale_k),	
	.fifo_scale_rden    (fifo_rden),
	.pixel_data         ({pixel_data[15:11],3'b0}),
	.sram_data_out      (data_out_r),
	.data_valid         (data_valid),
	.fifo_scale_rdempty (fifo_empty_r)
);      

//��ɫ��������ģ��      
 vin_scale_down u_vin_scale_down_g(
	.pixel_clk          (pixel_clk),
	.sram_clk           (sram_clk),
	.sys_rst_n          (sys_rst_n),	
	.hs                 (hs),
	.vs                 (vs),
	.de                 (de),
    .s_width            (s_width),
    .s_height           (s_height),
    .t_width            (t_width),
    .t_height           (t_height),
	.h_scale_k          (h_scale_k),
	.v_scale_k          (v_scale_k),		
	.fifo_scale_rden    (fifo_rden),	
	.pixel_data         ({pixel_data[10:5],2'b0}),
	.sram_data_out      (data_out_g),
	.data_valid         (),
    .fifo_scale_rdempty (fifo_empty_g)
);     

//��ɫ��������ģ�� 
 vin_scale_down u_vin_scale_down_b(
	.pixel_clk          (pixel_clk),
	.sram_clk           (sram_clk),	
	.sys_rst_n          (sys_rst_n),	
	.hs                 (hs),
	.vs                 (vs),
	.de                 (de),
    .s_width            (s_width),
    .s_height           (s_height),
    .t_width            (t_width),
    .t_height           (t_height),
	.h_scale_k          (h_scale_k),
	.v_scale_k          (v_scale_k),	
	.fifo_scale_rden    (fifo_rden),		
	.pixel_data         ({pixel_data[4:0],3'b0}),
	.sram_data_out      (data_out_b),
	.data_valid         (),
	.fifo_scale_rdempty (fifo_empty_b)
);   
 
endmodule
